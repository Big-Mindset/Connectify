<svg width="76" height="53" viewBox="0 0 76 53" fill="none" xmlns="http://www.w3.org/2000/svg">
<path d="M62.5848 5.27246C62.9991 5.6535 63.0174 6.30117 62.6253 6.70499L23.6947 46.8045L17.2072 40.8366L56.1753 0.698451C56.5527 0.30971 57.1711 0.292242 57.5698 0.659058L62.5848 5.27246Z" fill="#D9D9D9"/>
<path d="M4.8066 26.935C5.17362 26.5223 5.8057 26.4852 6.21839 26.8522L25.8516 44.3121L21.045 49.717C20.678 50.1297 20.0459 50.1668 19.6332 49.7998L0.747246 33.0044C0.334549 32.6374 0.297516 32.0053 0.66453 31.5926L4.8066 26.935Z" fill="#D9D9D9"/>
<path d="M70.1373 6.87803C70.5304 6.49016 71.1636 6.49445 71.5514 6.88761L75.2235 10.6097C75.6113 11.0029 75.607 11.636 75.2139 12.0239L39.0884 47.6635L34.0117 42.5177L70.1373 6.87803Z" fill="#D9D9D9"/>
<path d="M25.6835 44.7419C25.4853 44.5497 25.4805 44.2331 25.6728 44.0349L30.1423 39.427C30.3345 39.2287 30.6511 39.2239 30.8493 39.4162L39.2154 47.5309L34.7459 52.1389C34.3614 52.5353 33.7283 52.545 33.3318 52.1604L25.6835 44.7419Z" fill="#D9D9D9"/>
</svg>
