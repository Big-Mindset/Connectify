<svg width="63" height="51" viewBox="0 0 63 51" fill="none" xmlns="http://www.w3.org/2000/svg">
<path d="M62.5849 5.27245C62.9991 5.65349 63.0174 6.30117 62.6253 6.70498L23.6947 46.8045L17.2072 40.8366L56.1753 0.698443C56.5527 0.309703 57.1711 0.292234 57.5698 0.659051L62.5849 5.27245Z" fill="#D9D9D9"/>
<path d="M4.80661 26.9349C5.17362 26.5222 5.8057 26.4852 6.2184 26.8522L25.8516 44.3121L21.045 49.717C20.678 50.1297 20.0459 50.1668 19.6332 49.7998L0.747254 33.0044C0.334556 32.6374 0.297524 32.0053 0.664537 31.5926L4.80661 26.9349Z" fill="#D9D9D9"/>
</svg>
